* Truth-table DC sweep for TNOR

.include '../models/sky130_models.spice'
.include '../cells/sti.spice'
.include '../cells/tmax.spice'
.include '../cells/tnor.spice'

.param VDD_NOM=1.8

VDD vdd 0 DC VDD_NOM
VSS vss 0 DC 0

VA a 0 DC 0
VB b 0 DC 0

XTNOR a b y vdd vss TNOR

.dc VA 0 1.8 0.9 VB 0 1.8 0.9

.control
  run
  set filetype=ascii
  wrdata ../results/tnor_dc.csv V(a) V(b) V(y)
  quit
.endc

.end
