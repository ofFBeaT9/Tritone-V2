// BTISA Instruction Decoder
// Decodes 9-trit instructions for Balanced Ternary CPU
//
// Instruction format (9 trits):
//   [8:6] Opcode  (3 trits)
//   [5:4] Rd      (2 trits)
//   [3:2] Rs1     (2 trits)
//   [1:0] Rs2/Imm (2 trits)

`include "ternary_defs.vh"

module btisa_decoder (
  input  wire [17:0] instruction,  // 9 trits = 18 bits

  // Decoded fields
  output wire [5:0]  opcode,       // 3 trits = 6 bits
  output wire [3:0]  rd,           // 2 trits = 4 bits
  output wire [3:0]  rs1,          // 2 trits = 4 bits
  output wire [3:0]  rs2_imm,      // 2 trits = 4 bits

  // Control signals
  output reg         reg_write,
  output reg         mem_read,
  output reg         mem_write,
  output reg         branch,
  output reg         jump,
  output reg         alu_src,
  output reg  [2:0]  alu_op,
  output reg         halt
);

  // Extract instruction fields
  assign opcode  = instruction[17:12];  // Trits 8:6
  assign rd      = instruction[11:8];   // Trits 5:4
  assign rs1     = instruction[7:4];    // Trits 3:2
  assign rs2_imm = instruction[3:0];    // Trits 1:0

  // Opcode comparison helpers - compare 3 trits (6 bits)
  wire op_is_add  = (opcode == {`T_ZERO, `T_ZERO, `T_ZERO});       // 000
  wire op_is_sub  = (opcode == {`T_ZERO, `T_ZERO, `T_POS_ONE});    // 00+
  wire op_is_neg  = (opcode == {`T_ZERO, `T_ZERO, `T_NEG_ONE});    // 00-
  wire op_is_mul  = (opcode == {`T_ZERO, `T_POS_ONE, `T_ZERO});    // 0+0
  wire op_is_shl  = (opcode == {`T_ZERO, `T_POS_ONE, `T_POS_ONE}); // 0++
  wire op_is_shr  = (opcode == {`T_ZERO, `T_POS_ONE, `T_NEG_ONE}); // 0+-
  wire op_is_addi = (opcode == {`T_ZERO, `T_NEG_ONE, `T_ZERO});    // 0-0

  wire op_is_beq  = (opcode == {`T_ZERO, `T_NEG_ONE, `T_ZERO});    // 0-0
  wire op_is_bne  = (opcode == {`T_ZERO, `T_NEG_ONE, `T_POS_ONE}); // 0-+
  wire op_is_blt  = (opcode == {`T_ZERO, `T_NEG_ONE, `T_NEG_ONE}); // 0--

  wire op_is_min  = (opcode == {`T_POS_ONE, `T_ZERO, `T_ZERO});    // +00
  wire op_is_max  = (opcode == {`T_POS_ONE, `T_ZERO, `T_POS_ONE}); // +0+
  wire op_is_xor  = (opcode == {`T_POS_ONE, `T_ZERO, `T_NEG_ONE}); // +0-
  wire op_is_inv  = (opcode == {`T_POS_ONE, `T_POS_ONE, `T_ZERO}); // ++0
  wire op_is_pti  = (opcode == {`T_POS_ONE, `T_POS_ONE, `T_POS_ONE}); // +++
  wire op_is_nti  = (opcode == {`T_POS_ONE, `T_POS_ONE, `T_NEG_ONE}); // ++-

  wire op_is_jal  = (opcode == {`T_POS_ONE, `T_NEG_ONE, `T_ZERO});    // +-0
  wire op_is_jalr = (opcode == {`T_POS_ONE, `T_NEG_ONE, `T_POS_ONE}); // +-+
  wire op_is_jr   = (opcode == {`T_POS_ONE, `T_NEG_ONE, `T_NEG_ONE}); // +--

  wire op_is_ld   = (opcode == {`T_NEG_ONE, `T_ZERO, `T_ZERO});       // -00
  wire op_is_st   = (opcode == {`T_NEG_ONE, `T_ZERO, `T_POS_ONE});    // -0+
  wire op_is_ldt  = (opcode == {`T_NEG_ONE, `T_ZERO, `T_NEG_ONE});    // -0-
  wire op_is_stt  = (opcode == {`T_NEG_ONE, `T_POS_ONE, `T_ZERO});    // -+0
  wire op_is_lui  = (opcode == {`T_NEG_ONE, `T_POS_ONE, `T_POS_ONE}); // -++

  wire op_is_nop  = (opcode == {`T_NEG_ONE, `T_NEG_ONE, `T_ZERO});    // --0
  wire op_is_ecall= (opcode == {`T_NEG_ONE, `T_NEG_ONE, `T_NEG_ONE}); // ---
  wire op_is_halt = (opcode == {`T_NEG_ONE, `T_NEG_ONE, `T_POS_ONE}); // --+

  // Group classifications
  wire is_arithmetic = op_is_add | op_is_sub | op_is_neg | op_is_mul | op_is_shl | op_is_shr;
  wire is_logic      = op_is_min | op_is_max | op_is_xor | op_is_inv | op_is_pti | op_is_nti;
  wire is_branch     = op_is_beq | op_is_bne | op_is_blt;
  wire is_jump       = op_is_jal | op_is_jalr | op_is_jr;
  wire is_memory     = op_is_ld | op_is_st | op_is_ldt | op_is_stt | op_is_lui;

  // Decode control signals
  always @(*) begin
    // Defaults
    reg_write = 1'b0;
    mem_read  = 1'b0;
    mem_write = 1'b0;
    branch    = 1'b0;
    jump      = 1'b0;
    alu_src   = 1'b0;
    alu_op    = 3'b000;
    halt      = 1'b0;

    // Arithmetic operations
    if (is_arithmetic) begin
      reg_write = 1'b1;
      alu_src   = 1'b1;
      if (op_is_add)      alu_op = 3'b000;
      else if (op_is_sub) alu_op = 3'b001;
      else if (op_is_neg) alu_op = 3'b010;
      else if (op_is_mul) alu_op = 3'b000;
      else if (op_is_shl) alu_op = 3'b101;
      else if (op_is_shr) alu_op = 3'b110;
      else                alu_op = 3'b000;
    end

    // Logic operations
    if (is_logic) begin
      reg_write = 1'b1;
      if (op_is_min)      alu_op = 3'b011;
      else if (op_is_max) alu_op = 3'b100;
      else if (op_is_xor) alu_op = 3'b000;
      else if (op_is_inv) alu_op = 3'b010;
      else if (op_is_pti) alu_op = 3'b010;
      else if (op_is_nti) alu_op = 3'b010;
      else                alu_op = 3'b011;
    end

    // Branch operations
    if (is_branch) begin
      branch = 1'b1;
      alu_op = 3'b001;
    end

    // Jump operations
    if (is_jump) begin
      jump = 1'b1;
      if (op_is_jal || op_is_jalr) begin
        reg_write = 1'b1;
      end
      alu_op  = 3'b000;
      alu_src = 1'b1;
    end

    // Memory operations
    if (op_is_ld || op_is_ldt) begin
      reg_write = 1'b1;
      mem_read  = 1'b1;
      alu_src   = 1'b1;
      alu_op    = 3'b000;
    end

    if (op_is_st || op_is_stt) begin
      mem_write = 1'b1;
      alu_src   = 1'b1;
      alu_op    = 3'b000;
    end

    if (op_is_lui) begin
      reg_write = 1'b1;
      alu_src   = 1'b1;
    end

    // System operations
    if (op_is_halt) begin
      halt = 1'b1;
    end
  end

endmodule
