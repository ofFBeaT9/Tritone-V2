* ============================================================================
* Testbench for 3-Rail STI
* ============================================================================

.include '../cells/sti_3rail.spice'

* Power supplies
VDD  vdd  0 DC 1.8
VMID vmid 0 DC 0.9
VSS  vss  0 DC 0

* DC sweep input
VIN_DC in_dc 0 DC 0

* Transient input - test all transitions
VIN_TR in_tr 0 PWL(0n 0 20n 0 30n 0.9 50n 0.9 60n 1.8 80n 1.8 90n 0.9 110n 0.9 120n 0)

* Device under test - DC
XSTI_DC in_dc out_dc vdd vmid vss STI_3RAIL
CL_DC out_dc 0 20f

* Device under test - Transient
XSTI_TR in_tr out_tr vdd vmid vss STI_3RAIL
CL_TR out_tr 0 20f

* DC sweep analysis
.dc VIN_DC 0 1.8 0.01

* Transient analysis
.tran 0.1n 120n

* Measurements
.meas DC vout_at_0 FIND V(out_dc) AT=0
.meas DC vout_at_mid FIND V(out_dc) AT=0.9
.meas DC vout_at_high FIND V(out_dc) AT=1.8

.control
run

echo ""
echo "=============================================="
echo "3-Rail STI Test Results"
echo "=============================================="
echo ""

set filetype=ascii

* DC transfer curve
setplot dc1
echo "DC Transfer Characteristic:"
echo "  Vin=0V    -> Vout should be ~1.8V"
echo "  Vin=0.9V  -> Vout should be ~0.9V"
echo "  Vin=1.8V  -> Vout should be ~0V"
echo ""

* Save DC results
wrdata ../results/sti_3rail_dc.csv V(out_dc)

* Transient results
setplot tran1
echo "Transient test completed"
wrdata ../results/sti_3rail_tran.csv V(in_tr) V(out_tr)

echo ""
echo "Results saved to ../results/"
echo ""

quit

.endc

.end
