* ============================================================================
* MONTE CARLO ANALYSIS FOR STI
* ============================================================================
* GT-LOGIC Ternary CMOS Cell Library
* Process Variation Analysis for Standard Ternary Inverter
*
* Tests:
*   1. Vth variation impact on output levels
*   2. Sizing mismatch effects
*   3. Statistical distribution of mid-level voltage
*   4. 3-sigma yield estimation
* ============================================================================

.include '../models/sky130_models.spice'
.include '../cells/sti.spice'

* ============================================================================
* POWER SUPPLIES (2-rail)
* ============================================================================
VDD vdd 0 DC 1.8
VSS vss 0 DC 0

* ============================================================================
* TEST INPUT AT MID-LEVEL (Most sensitive point)
* ============================================================================
VIN in 0 DC 0.9

* ============================================================================
* DEVICE UNDER TEST
* ============================================================================
XSTI in out vdd vss STI

* Load capacitance
CL out 0 20f

* ============================================================================
* PROCESS VARIATION PARAMETERS
* ============================================================================
* Typical 3-sigma variations for 130nm technology:
*   Vth: ±30mV (σ = 10mV)
*   Tox: ±5% (σ = 1.67%)
*   W/L: ±5% (σ = 1.67%)

.param vth_nom = 0.42
.param vth_sigma = 0.010
.param tox_nom = 4.15e-9
.param tox_sigma_pct = 0.0167
.param wl_sigma_pct = 0.0167

* ============================================================================
* DC ANALYSIS
* ============================================================================
.dc VIN 0 1.8 0.01

* Key measurements
.meas DC vout_at_0 FIND V(out) AT=0
.meas DC vout_at_mid FIND V(out) AT=0.9
.meas DC vout_at_high FIND V(out) AT=1.8
.meas DC switching_threshold WHEN V(out)=0.9 CROSS=1

* ============================================================================
* SIMULATION CONTROL WITH MONTE CARLO
* ============================================================================
.control
    * Run nominal DC sweep first
    run
    
    echo ""
    echo "============================================================"
    echo "STI MONTE CARLO PROCESS VARIATION ANALYSIS"
    echo "============================================================"
    echo ""
    
    * Store nominal results
    setplot dc1
    let vout_nom = V(out)
    
    echo "=== Nominal Results ==="
    echo "Vout at Vin=0V:   should be ~1.8V"
    echo "Vout at Vin=0.9V: should be ~0.9V"
    echo "Vout at Vin=1.8V: should be ~0V"
    echo ""
    
    * Plot nominal transfer curve
    plot vout_nom vs V(in) title 'STI Nominal DC Transfer Curve'
    
    echo ""
    echo "=== Process Variation Analysis ==="
    echo ""
    echo "For full Monte Carlo, run with ngspice -b with .param variations"
    echo "This requires updating model parameters in a loop"
    echo ""
    echo "Key metrics to track:"
    echo "  - Vout at Vin=0.9V: Target 0.9V ± 50mV"
    echo "  - Switching threshold: Target 0.9V ± 100mV"
    echo "  - Gain at mid-point: Higher is better"
    echo ""
    
    * Calculate gain at mid-point (slope of transfer curve)
    let deriv_vout = deriv(vout_nom)
    let gain_at_mid = -deriv_vout[90]
    echo "Gain at Vin=0.9V (nominal): " gain_at_mid
    echo ""
    
    * Noise margin calculation
    * NML = VIL - VOL (low noise margin)
    * NMH = VOH - VIH (high noise margin)
    * For ternary, we have additional margins for intermediate level
    
    echo "=== Noise Margins ==="
    let vol = vout_nom[180]
    let voh = vout_nom[0]
    let vom = vout_nom[90]
    
    echo "VOL (Vout at Vin=1.8V): " vol
    echo "VOH (Vout at Vin=0V): " voh
    echo "VOM (Vout at Vin=0.9V): " vom
    echo ""
    
    * Ternary noise margins (simplified)
    * NM_low = (0.45V threshold) - VOL
    * NM_high = VOH - (1.35V threshold)
    * NM_mid = min(VOM - 0.45V, 1.35V - VOM)
    
    let nm_low = 0.45 - vol
    let nm_high = voh - 1.35
    let nm_mid_lo = vom - 0.45
    let nm_mid_hi = 1.35 - vom
    
    echo "Ternary Noise Margins:"
    echo "  NM_low:  " nm_low " V"
    echo "  NM_high: " nm_high " V"
    echo "  NM_mid (lower boundary): " nm_mid_lo " V"
    echo "  NM_mid (upper boundary): " nm_mid_hi " V"
    echo ""
    
    echo "=== Verification Criteria ==="
    echo "  ✓ Vout at Vin=0.9V within [0.85V, 0.95V]: PASS if VOM in range"
    echo "  ✓ All noise margins > 100mV: PASS if NM > 0.1V"
    echo "  ✓ Gain at mid-point > 1: PASS if gain > 1"
    echo ""
    
    * Save results
    wrdata ../results/sti_monte_carlo.csv vout_nom
    
    echo "Nominal curve saved to ../results/sti_monte_carlo.csv"
    echo ""
    echo "For production Monte Carlo analysis:"
    echo "  1. Use .param statements with GAUSS() function"
    echo "  2. Run 1000+ iterations"
    echo "  3. Analyze distribution of Vout at Vin=0.9V"
    echo "  4. Calculate yield for ±50mV specification"
    echo ""
    quit
.endc

.end
